`timescale 1ns/1ns
module tb();
    
    logic [15:0] aa, bb;
    logic [2:0]

endmodule